-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0b95",
     9 => x"88080b0b",
    10 => x"0b958c08",
    11 => x"0b0b0b95",
    12 => x"90080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"95900c0b",
    16 => x"0b0b958c",
    17 => x"0c0b0b0b",
    18 => x"95880c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b94d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"95887099",
    57 => x"e0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"dc050d83",
    63 => x"a82d840b",
    64 => x"ec0c8b82",
    65 => x"2d958808",
    66 => x"53958808",
    67 => x"802e818f",
    68 => x"38850bec",
    69 => x"0c94e452",
    70 => x"95985191",
    71 => x"aa2d9588",
    72 => x"08802e80",
    73 => x"f438959c",
    74 => x"0870f80c",
    75 => x"ff115457",
    76 => x"72802e88",
    77 => x"3872812a",
    78 => x"5382b004",
    79 => x"80772580",
    80 => x"d83895a8",
    81 => x"52959851",
    82 => x"93e02d95",
    83 => x"8808802e",
    84 => x"b83895a8",
    85 => x"5983fc58",
    86 => x"78708405",
    87 => x"5a087081",
    88 => x"ff067188",
    89 => x"2a7081ff",
    90 => x"0673902a",
    91 => x"7081ff06",
    92 => x"75982ae8",
    93 => x"0ce80c58",
    94 => x"e80c57e8",
    95 => x"0cfc1959",
    96 => x"53778025",
    97 => x"d338838c",
    98 => x"04848057",
    99 => x"95985193",
   100 => x"b32dfc80",
   101 => x"175782bc",
   102 => x"04840bec",
   103 => x"0c805372",
   104 => x"95880c02",
   105 => x"a4050d04",
   106 => x"810bffb0",
   107 => x"0c0402f4",
   108 => x"050dd452",
   109 => x"81ff720c",
   110 => x"71085381",
   111 => x"ff720c72",
   112 => x"882b83fe",
   113 => x"80067208",
   114 => x"7081ff06",
   115 => x"51525381",
   116 => x"ff720c72",
   117 => x"7107882b",
   118 => x"72087081",
   119 => x"ff065152",
   120 => x"5381ff72",
   121 => x"0c727107",
   122 => x"882b7208",
   123 => x"7081ff06",
   124 => x"72079588",
   125 => x"0c525302",
   126 => x"8c050d04",
   127 => x"02f4050d",
   128 => x"74767181",
   129 => x"ff06d40c",
   130 => x"535395a4",
   131 => x"08853871",
   132 => x"892b5271",
   133 => x"982ad40c",
   134 => x"71902a70",
   135 => x"81ff06d4",
   136 => x"0c517188",
   137 => x"2a7081ff",
   138 => x"06d40c51",
   139 => x"7181ff06",
   140 => x"d40c7290",
   141 => x"2a7081ff",
   142 => x"06d40c51",
   143 => x"d4087081",
   144 => x"ff065151",
   145 => x"82b8bf52",
   146 => x"7081ff2e",
   147 => x"09810694",
   148 => x"3881ff0b",
   149 => x"d40cd408",
   150 => x"7081ff06",
   151 => x"ff145451",
   152 => x"5171e538",
   153 => x"7095880c",
   154 => x"028c050d",
   155 => x"0402fc05",
   156 => x"0d81c751",
   157 => x"81ff0bd4",
   158 => x"0cff1151",
   159 => x"708025f4",
   160 => x"38028405",
   161 => x"0d0402f4",
   162 => x"050d81ff",
   163 => x"0bd40c93",
   164 => x"53805287",
   165 => x"fc80c151",
   166 => x"83fc2d95",
   167 => x"88088b38",
   168 => x"81ff0bd4",
   169 => x"0c815385",
   170 => x"b30484ed",
   171 => x"2dff1353",
   172 => x"72df3872",
   173 => x"95880c02",
   174 => x"8c050d04",
   175 => x"02ec050d",
   176 => x"810b95a4",
   177 => x"0c8454d0",
   178 => x"08708f2a",
   179 => x"70810651",
   180 => x"515372f3",
   181 => x"3872d00c",
   182 => x"84ed2dd0",
   183 => x"08708f2a",
   184 => x"70810651",
   185 => x"515372f3",
   186 => x"38810bd0",
   187 => x"0cb15380",
   188 => x"5284d480",
   189 => x"c05183fc",
   190 => x"2d958808",
   191 => x"812e9338",
   192 => x"72822ebd",
   193 => x"38ff1353",
   194 => x"72e538ff",
   195 => x"145473ff",
   196 => x"b63884ed",
   197 => x"2d83aa52",
   198 => x"849c80c8",
   199 => x"5183fc2d",
   200 => x"95880881",
   201 => x"2e098106",
   202 => x"923883ae",
   203 => x"2d958808",
   204 => x"83ffff06",
   205 => x"537283aa",
   206 => x"2e913885",
   207 => x"862d86c6",
   208 => x"04805388",
   209 => x"94048054",
   210 => x"87e60481",
   211 => x"ff0bd40c",
   212 => x"b15484ed",
   213 => x"2d8fcf53",
   214 => x"805287fc",
   215 => x"80f75183",
   216 => x"fc2d9588",
   217 => x"08559588",
   218 => x"08812e09",
   219 => x"81069b38",
   220 => x"81ff0bd4",
   221 => x"0c820a52",
   222 => x"849c80e9",
   223 => x"5183fc2d",
   224 => x"95880880",
   225 => x"2e8d3884",
   226 => x"ed2dff13",
   227 => x"5372c938",
   228 => x"87d90481",
   229 => x"ff0bd40c",
   230 => x"95880852",
   231 => x"87fc80fa",
   232 => x"5183fc2d",
   233 => x"958808b1",
   234 => x"3881ff0b",
   235 => x"d40cd408",
   236 => x"5381ff0b",
   237 => x"d40c81ff",
   238 => x"0bd40c81",
   239 => x"ff0bd40c",
   240 => x"81ff0bd4",
   241 => x"0c72862a",
   242 => x"70810676",
   243 => x"56515372",
   244 => x"95389588",
   245 => x"085487e6",
   246 => x"0473822e",
   247 => x"fee838ff",
   248 => x"145473fe",
   249 => x"ed387395",
   250 => x"a40c738b",
   251 => x"38815287",
   252 => x"fc80d051",
   253 => x"83fc2d81",
   254 => x"ff0bd40c",
   255 => x"d008708f",
   256 => x"2a708106",
   257 => x"51515372",
   258 => x"f33872d0",
   259 => x"0c81ff0b",
   260 => x"d40c8153",
   261 => x"7295880c",
   262 => x"0294050d",
   263 => x"0402e805",
   264 => x"0d785580",
   265 => x"5681ff0b",
   266 => x"d40cd008",
   267 => x"708f2a70",
   268 => x"81065151",
   269 => x"5372f338",
   270 => x"82810bd0",
   271 => x"0c81ff0b",
   272 => x"d40c7752",
   273 => x"87fc80d1",
   274 => x"5183fc2d",
   275 => x"95880880",
   276 => x"d93880db",
   277 => x"c6df5481",
   278 => x"ff0bd40c",
   279 => x"d4087081",
   280 => x"ff065153",
   281 => x"7281fe2e",
   282 => x"0981069d",
   283 => x"3880ff53",
   284 => x"83ae2d95",
   285 => x"88087570",
   286 => x"8405570c",
   287 => x"ff135372",
   288 => x"8025ed38",
   289 => x"8156898f",
   290 => x"04ff1454",
   291 => x"73c93881",
   292 => x"ff0bd40c",
   293 => x"81ff0bd4",
   294 => x"0cd00870",
   295 => x"8f2a7081",
   296 => x"06515153",
   297 => x"72f33872",
   298 => x"d00c7595",
   299 => x"880c0298",
   300 => x"050d0402",
   301 => x"e8050d77",
   302 => x"797b5855",
   303 => x"55805372",
   304 => x"7625a338",
   305 => x"74708105",
   306 => x"5680f52d",
   307 => x"74708105",
   308 => x"5680f52d",
   309 => x"52527171",
   310 => x"2e863881",
   311 => x"5189e804",
   312 => x"81135389",
   313 => x"bf048051",
   314 => x"7095880c",
   315 => x"0298050d",
   316 => x"0402ec05",
   317 => x"0d765574",
   318 => x"802ebb38",
   319 => x"9a1580e0",
   320 => x"2d5194b6",
   321 => x"2d958808",
   322 => x"95880899",
   323 => x"d40c9588",
   324 => x"08545499",
   325 => x"b008802e",
   326 => x"99389415",
   327 => x"80e02d51",
   328 => x"94b62d95",
   329 => x"8808902b",
   330 => x"83fff00a",
   331 => x"06707507",
   332 => x"51537299",
   333 => x"d40c99d4",
   334 => x"08537280",
   335 => x"2e993899",
   336 => x"a808fe14",
   337 => x"712999bc",
   338 => x"080599d8",
   339 => x"0c70842b",
   340 => x"99b40c54",
   341 => x"8afd0499",
   342 => x"c00899d4",
   343 => x"0c99c408",
   344 => x"99d80c99",
   345 => x"b008802e",
   346 => x"8a3899a8",
   347 => x"08842b53",
   348 => x"8af90499",
   349 => x"c808842b",
   350 => x"537299b4",
   351 => x"0c029405",
   352 => x"0d0402d8",
   353 => x"050d800b",
   354 => x"99b00c84",
   355 => x"5485bc2d",
   356 => x"95880880",
   357 => x"2e953895",
   358 => x"a8528051",
   359 => x"889d2d95",
   360 => x"8808802e",
   361 => x"8638fe54",
   362 => x"8bb304ff",
   363 => x"14547380",
   364 => x"24db3873",
   365 => x"5573802e",
   366 => x"84f93880",
   367 => x"56810b99",
   368 => x"dc0c8853",
   369 => x"94f05295",
   370 => x"de5189b3",
   371 => x"2d958808",
   372 => x"762e0981",
   373 => x"06873895",
   374 => x"880899dc",
   375 => x"0c885394",
   376 => x"fc5295fa",
   377 => x"5189b32d",
   378 => x"95880887",
   379 => x"38958808",
   380 => x"99dc0c99",
   381 => x"dc08802e",
   382 => x"80f63898",
   383 => x"ee0b80f5",
   384 => x"2d98ef0b",
   385 => x"80f52d71",
   386 => x"982b7190",
   387 => x"2b0798f0",
   388 => x"0b80f52d",
   389 => x"70882b72",
   390 => x"0798f10b",
   391 => x"80f52d71",
   392 => x"0799a60b",
   393 => x"80f52d99",
   394 => x"a70b80f5",
   395 => x"2d71882b",
   396 => x"07535f54",
   397 => x"525a5657",
   398 => x"557381ab",
   399 => x"aa2e0981",
   400 => x"068d3875",
   401 => x"5194862d",
   402 => x"95880856",
   403 => x"8cdc0480",
   404 => x"557382d4",
   405 => x"d52e0981",
   406 => x"0683d838",
   407 => x"95a85275",
   408 => x"51889d2d",
   409 => x"95880855",
   410 => x"95880880",
   411 => x"2e83c438",
   412 => x"885394fc",
   413 => x"5295fa51",
   414 => x"89b32d95",
   415 => x"88088938",
   416 => x"810b99b0",
   417 => x"0c8da004",
   418 => x"885394f0",
   419 => x"5295de51",
   420 => x"89b32d80",
   421 => x"55958808",
   422 => x"752e0981",
   423 => x"06839438",
   424 => x"99a60b80",
   425 => x"f52d5473",
   426 => x"80d52e09",
   427 => x"810680ca",
   428 => x"3899a70b",
   429 => x"80f52d54",
   430 => x"7381aa2e",
   431 => x"098106ba",
   432 => x"38800b95",
   433 => x"a80b80f5",
   434 => x"2d565474",
   435 => x"81e92e83",
   436 => x"38815474",
   437 => x"81eb2e8c",
   438 => x"38805573",
   439 => x"752e0981",
   440 => x"0682d038",
   441 => x"95b30b80",
   442 => x"f52d5574",
   443 => x"8d3895b4",
   444 => x"0b80f52d",
   445 => x"5473822e",
   446 => x"86388055",
   447 => x"90b30495",
   448 => x"b50b80f5",
   449 => x"2d7099a8",
   450 => x"0cff0599",
   451 => x"ac0c95b6",
   452 => x"0b80f52d",
   453 => x"95b70b80",
   454 => x"f52d5876",
   455 => x"05778280",
   456 => x"29057099",
   457 => x"b80c95b8",
   458 => x"0b80f52d",
   459 => x"7099cc0c",
   460 => x"99b00859",
   461 => x"57587680",
   462 => x"2e81a338",
   463 => x"885394fc",
   464 => x"5295fa51",
   465 => x"89b32d95",
   466 => x"880881e7",
   467 => x"3899a808",
   468 => x"70842b99",
   469 => x"b40c7099",
   470 => x"c80c95cd",
   471 => x"0b80f52d",
   472 => x"95cc0b80",
   473 => x"f52d7182",
   474 => x"80290595",
   475 => x"ce0b80f5",
   476 => x"2d708480",
   477 => x"80291295",
   478 => x"cf0b80f5",
   479 => x"2d708180",
   480 => x"0a291270",
   481 => x"99d00c99",
   482 => x"cc087129",
   483 => x"99b80805",
   484 => x"7099bc0c",
   485 => x"95d50b80",
   486 => x"f52d95d4",
   487 => x"0b80f52d",
   488 => x"71828029",
   489 => x"0595d60b",
   490 => x"80f52d70",
   491 => x"84808029",
   492 => x"1295d70b",
   493 => x"80f52d70",
   494 => x"982b81f0",
   495 => x"0a067205",
   496 => x"7099c00c",
   497 => x"fe117e29",
   498 => x"770599c4",
   499 => x"0c525952",
   500 => x"43545e51",
   501 => x"5259525d",
   502 => x"57595790",
   503 => x"ac0495ba",
   504 => x"0b80f52d",
   505 => x"95b90b80",
   506 => x"f52d7182",
   507 => x"80290570",
   508 => x"99b40c70",
   509 => x"a02983ff",
   510 => x"0570892a",
   511 => x"7099c80c",
   512 => x"95bf0b80",
   513 => x"f52d95be",
   514 => x"0b80f52d",
   515 => x"71828029",
   516 => x"057099d0",
   517 => x"0c7b7129",
   518 => x"1e7099c4",
   519 => x"0c7d99c0",
   520 => x"0c730599",
   521 => x"bc0c555e",
   522 => x"51515555",
   523 => x"805189f1",
   524 => x"2d815574",
   525 => x"95880c02",
   526 => x"a8050d04",
   527 => x"02ec050d",
   528 => x"7670872c",
   529 => x"7180ff06",
   530 => x"55565499",
   531 => x"b0088a38",
   532 => x"73882c74",
   533 => x"81ff0654",
   534 => x"5595a852",
   535 => x"99b80815",
   536 => x"51889d2d",
   537 => x"95880854",
   538 => x"95880880",
   539 => x"2eb33899",
   540 => x"b008802e",
   541 => x"98387284",
   542 => x"2995a805",
   543 => x"70085253",
   544 => x"94862d95",
   545 => x"8808f00a",
   546 => x"0653919f",
   547 => x"04721095",
   548 => x"a8057080",
   549 => x"e02d5253",
   550 => x"94b62d95",
   551 => x"88085372",
   552 => x"54739588",
   553 => x"0c029405",
   554 => x"0d0402cc",
   555 => x"050d7e60",
   556 => x"5e5a800b",
   557 => x"99d40899",
   558 => x"d808595c",
   559 => x"56805899",
   560 => x"b408782e",
   561 => x"81ae3877",
   562 => x"8f06a017",
   563 => x"5754738f",
   564 => x"3895a852",
   565 => x"76518117",
   566 => x"57889d2d",
   567 => x"95a85680",
   568 => x"7680f52d",
   569 => x"56547474",
   570 => x"2e833881",
   571 => x"547481e5",
   572 => x"2e80f638",
   573 => x"81707506",
   574 => x"555c7380",
   575 => x"2e80ea38",
   576 => x"8b1680f5",
   577 => x"2d980659",
   578 => x"7880de38",
   579 => x"8b537c52",
   580 => x"755189b3",
   581 => x"2d958808",
   582 => x"80cf389c",
   583 => x"16085194",
   584 => x"862d9588",
   585 => x"08841b0c",
   586 => x"9a1680e0",
   587 => x"2d5194b6",
   588 => x"2d958808",
   589 => x"95880888",
   590 => x"1c0c9588",
   591 => x"08555599",
   592 => x"b008802e",
   593 => x"98389416",
   594 => x"80e02d51",
   595 => x"94b62d95",
   596 => x"8808902b",
   597 => x"83fff00a",
   598 => x"06701651",
   599 => x"5473881b",
   600 => x"0c787a0c",
   601 => x"7b5493aa",
   602 => x"04811858",
   603 => x"99b40878",
   604 => x"26fed438",
   605 => x"99b00880",
   606 => x"2eae387a",
   607 => x"5190bc2d",
   608 => x"95880895",
   609 => x"880880ff",
   610 => x"fffff806",
   611 => x"555b7380",
   612 => x"fffffff8",
   613 => x"2e923895",
   614 => x"8808fe05",
   615 => x"99a80829",
   616 => x"99bc0805",
   617 => x"5791bd04",
   618 => x"80547395",
   619 => x"880c02b4",
   620 => x"050d0402",
   621 => x"f4050d74",
   622 => x"70088105",
   623 => x"710c7008",
   624 => x"99ac0806",
   625 => x"5353718e",
   626 => x"38881308",
   627 => x"5190bc2d",
   628 => x"95880888",
   629 => x"140c810b",
   630 => x"95880c02",
   631 => x"8c050d04",
   632 => x"02f0050d",
   633 => x"75881108",
   634 => x"fe0599a8",
   635 => x"082999bc",
   636 => x"08117208",
   637 => x"99ac0806",
   638 => x"05795553",
   639 => x"5454889d",
   640 => x"2d029005",
   641 => x"0d0402f4",
   642 => x"050d7470",
   643 => x"882a83fe",
   644 => x"80067072",
   645 => x"982a0772",
   646 => x"882b87fc",
   647 => x"80800673",
   648 => x"982b81f0",
   649 => x"0a067173",
   650 => x"07079588",
   651 => x"0c565153",
   652 => x"51028c05",
   653 => x"0d0402f8",
   654 => x"050d028e",
   655 => x"0580f52d",
   656 => x"74882b07",
   657 => x"7083ffff",
   658 => x"0695880c",
   659 => x"51028805",
   660 => x"0d040000",
   661 => x"00ffffff",
   662 => x"ff00ffff",
   663 => x"ffff00ff",
   664 => x"ffffff00",
   665 => x"53504543",
   666 => x"5452554d",
   667 => x"524f4d00",
   668 => x"46415431",
   669 => x"36202020",
   670 => x"00000000",
   671 => x"46415433",
   672 => x"32202020",
   673 => x"00202020",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

